module MI(
	// IN
	input[31:0] I,  // Endereco da instrucao
	
	// OUT
	output[31:0] ID // Instrucao
	
	);
	// TODO: Alterar o tamanho da memória de instrução
	
	reg[31:0] mem_i[300:0];  // Memoria de fato
	
	initial begin
		/*
		// Gcd
		mem_i[0] = 32'b00000000000000000000000000000000;
		mem_i[1] = 32'b00010111101000000010010101100000;
		mem_i[2] = 32'b00000111101111111111111111100011;
		mem_i[3] = 32'b00011011101111110000000000000000;
		mem_i[4] = 32'b00000111101111111111111111100011;
		mem_i[5] = 32'b00011011101111000000000000000000;
		mem_i[6] = 32'b00010011100111010000000000000000;
		mem_i[7] = 32'b00000111101111111111111111100011;
		mem_i[8] = 32'b00000111101111111111111111100011;
		mem_i[9] = 32'b00010001001111000000000000000000;
		mem_i[10] = 32'b00011101001000001111111111111111;
		mem_i[11] = 32'b00010111011000000000000000000000;
		mem_i[12] = 32'b01000011011000000000000000000000;
		mem_i[13] = 32'b00011111011000000000000000000000;
		mem_i[14] = 32'b00010001010110110000000000000000;
		mem_i[15] = 32'b00010001001010100000000000000000;
		mem_i[16] = 32'b00011011100010011111111111111111;
		mem_i[17] = 32'b00010001011111000000000000000000;
		mem_i[18] = 32'b00011101011000001111111111111110;
		mem_i[19] = 32'b00010111011000000000000000000000;
		mem_i[20] = 32'b01000011011000000000000000000000;
		mem_i[21] = 32'b00011111011000000000000000000000;
		mem_i[22] = 32'b00010001100110110000000000000000;
		mem_i[23] = 32'b00010001011011000000000000000000;
		mem_i[24] = 32'b00011011100010111111111111111110;
		mem_i[25] = 32'b00011011101010011111111111111111;
		mem_i[26] = 32'b00011011101010111111111111111110;
		mem_i[27] = 32'b00000111101111111111111111000011;
		mem_i[28] = 32'b00011011101010111111111111111100;
		mem_i[29] = 32'b00011011101010011111111111111101;
		mem_i[30] = 32'b00111000000000000000000000001010;
		mem_i[31] = 32'b00010001011111010000000000000000;
		mem_i[32] = 32'b00011101011000000000000000000000;
		mem_i[33] = 32'b00010001001111010000000000000000;
		mem_i[34] = 32'b00011101001000000000000000000001;
		mem_i[35] = 32'b00000111101000000000000001000011;
		mem_i[36] = 32'b00010001101110100000000000000000;
		mem_i[37] = 32'b00010111011000000000000000100000;
		mem_i[38] = 32'b00011011011011010000000000000000;
		mem_i[39] = 32'b01000111011000000000000000000000;
		mem_i[40] = 32'b11111100000000000000000000000000;
		mem_i[41] = 32'b00000111101111111111111111100011;
		mem_i[42] = 32'b00011011101111110000000000000000;
		mem_i[43] = 32'b00000111101111111111111111100011;
		mem_i[44] = 32'b00011011101111000000000000000000;
		mem_i[45] = 32'b00010011100111010000000000000000;
		mem_i[46] = 32'b00000111101111111111111111100011;
		mem_i[47] = 32'b00010000000111000000000000000000;
		mem_i[48] = 32'b00011100000000001111111111111111;
		mem_i[49] = 32'b00000111101111111111111111100011;
		mem_i[50] = 32'b00010000001111000000000000000000;
		mem_i[51] = 32'b00011100001000001111111111111110;
		mem_i[52] = 32'b00001100001000000000000000001001;
		mem_i[53] = 32'b00000111110000000000000000100011;
		mem_i[54] = 32'b00111100000000000000000000000010;
		mem_i[55] = 32'b00010011010000000000000000000000;
		mem_i[56] = 32'b00110100000000000000000000100000;
		mem_i[57] = 32'b00010000011111000000000000000000;
		mem_i[58] = 32'b00011100011000001111111111111110;
		mem_i[59] = 32'b00010000100111000000000000000000;
		mem_i[60] = 32'b00011100100000001111111111111111;
		mem_i[61] = 32'b00010011011001000000000000000000;
		mem_i[62] = 32'b00000111011000110000000000000110;
		mem_i[63] = 32'b00010000101110110000000000000000;
		mem_i[64] = 32'b00010011011001010000000000000000;
		mem_i[65] = 32'b00000111011000110000000000000101;
		mem_i[66] = 32'b00010000110110110000000000000000;
		mem_i[67] = 32'b00010011011001000000000000000000;
		mem_i[68] = 32'b00000111011001100000000000000010;
		mem_i[69] = 32'b00010000111110110000000000000000;
		mem_i[70] = 32'b00011011101000001111111111111111;
		mem_i[71] = 32'b00011011101000011111111111111110;
		mem_i[72] = 32'b00011011101000111111111111111101;
		mem_i[73] = 32'b00011011101001001111111111111100;
		mem_i[74] = 32'b00000111101111111111111110000011;
		mem_i[75] = 32'b00011011101001111111111111111100;
		mem_i[76] = 32'b00011011101000111111111111111101;
		mem_i[77] = 32'b00111000000000001111111111011011;
		mem_i[78] = 32'b00010000100111010000000000000000;
		mem_i[79] = 32'b00011100100000000000000000000000;
		mem_i[80] = 32'b00010000011111010000000000000000;
		mem_i[81] = 32'b00011100011000000000000000000001;
		mem_i[82] = 32'b00010000001111010000000000000000;
		mem_i[83] = 32'b00011100001000000000000000000010;
		mem_i[84] = 32'b00010000000111010000000000000000;
		mem_i[85] = 32'b00011100000000000000000000000011;
		mem_i[86] = 32'b00000111101000000000000010000011;
		mem_i[87] = 32'b00010001000110100000000000000000;
		mem_i[88] = 32'b00010011010010000000000000000000;
		mem_i[89] = 32'b00010011111111000000000000000000;
		mem_i[90] = 32'b00011111111000000000000000000001;
		mem_i[91] = 32'b00010011101111000000000000000000;
		mem_i[92] = 32'b00000111101000000000000001000011;
		mem_i[93] = 32'b00011111100000000000000000000000;
		mem_i[94] = 32'b00101011111000000000000000000000;
		*/
		/*
		//	Fatorial
		mem_i[0] = 32'b00000000000000000000000000000000;
		mem_i[1] = 32'b00010111101000000010010101100000;
		mem_i[2] = 32'b00000111101111111111111111100011;
		mem_i[3] = 32'b00011011101111110000000000000000;
		mem_i[4] = 32'b00000111101111111111111111100011;
		mem_i[5] = 32'b00011011101111000000000000000000;
		mem_i[6] = 32'b00010011100111010000000000000000;
		mem_i[7] = 32'b00000111101111111111111111100011;
		mem_i[8] = 32'b00010000110111000000000000000000;
		mem_i[9] = 32'b00011100110000001111111111111111;
		mem_i[10] = 32'b00010111011000000000000000000000;
		mem_i[11] = 32'b01000011011000000000000000000000;
		mem_i[12] = 32'b00011111011000000000000000000000;
		mem_i[13] = 32'b00010000111110110000000000000000;
		mem_i[14] = 32'b00010000110001110000000000000000;
		mem_i[15] = 32'b00011011100001101111111111111111;
		mem_i[16] = 32'b00011011101001101111111111111111;
		mem_i[17] = 32'b00000111101111111111111111100011;
		mem_i[18] = 32'b00011011101001101111111111111101;
		mem_i[19] = 32'b00111000000000000000000000001000;
		mem_i[20] = 32'b00010000110111010000000000000000;
		mem_i[21] = 32'b00011100110000000000000000000000;
		mem_i[22] = 32'b00000111101000000000000000100011;
		mem_i[23] = 32'b00010001000110100000000000000000;
		mem_i[24] = 32'b00010111011000000000000000100000;
		mem_i[25] = 32'b00011011011010000000000000000000;
		mem_i[26] = 32'b01000111011000000000000000000000;
		mem_i[27] = 32'b11111100000000000000000000000000;
		mem_i[28] = 32'b00000111101111111111111111100011;
		mem_i[29] = 32'b00011011101111110000000000000000;
		mem_i[30] = 32'b00000111101111111111111111100011;
		mem_i[31] = 32'b00011011101111000000000000000000;
		mem_i[32] = 32'b00010011100111010000000000000000;
		mem_i[33] = 32'b00000111101111111111111111100011;
		mem_i[34] = 32'b00010000000111000000000000000000;
		mem_i[35] = 32'b00011100000000001111111111111111;
		mem_i[36] = 32'b00001100000000000000000000001011;
		mem_i[37] = 32'b00000111110000000000000000100011;
		mem_i[38] = 32'b00111100000000000000000000000010;
		mem_i[39] = 32'b00010111010000000000000000100000;
		mem_i[40] = 32'b00110100000000000000000000010100;
		mem_i[41] = 32'b00010000010111000000000000000000;
		mem_i[42] = 32'b00011100010000001111111111111111;
		mem_i[43] = 32'b00010011011000100000000000000000;
		mem_i[44] = 32'b00000111011000000000000000100100;
		mem_i[45] = 32'b00010000011110110000000000000000;
		mem_i[46] = 32'b00011011101000001111111111111111;
		mem_i[47] = 32'b00011011101000101111111111111110;
		mem_i[48] = 32'b00000111101111111111111111000011;
		mem_i[49] = 32'b00011011101000111111111111111101;
		mem_i[50] = 32'b00111000000000001111111111101001;
		mem_i[51] = 32'b00010000010111010000000000000000;
		mem_i[52] = 32'b00011100010000000000000000000000;
		mem_i[53] = 32'b00010000000111010000000000000000;
		mem_i[54] = 32'b00011100000000000000000000000001;
		mem_i[55] = 32'b00000111101000000000000001000011;
		mem_i[56] = 32'b00010000100110100000000000000000;
		mem_i[57] = 32'b00010011011000100000000000000000;
		mem_i[58] = 32'b00000111011001000000000000000101;
		mem_i[59] = 32'b00010000101110110000000000000000;
		mem_i[60] = 32'b00010011010001010000000000000000;
		mem_i[61] = 32'b00010011111111000000000000000000;
		mem_i[62] = 32'b00011111111000000000000000000001;
		mem_i[63] = 32'b00010011101111000000000000000000;
		mem_i[64] = 32'b00000111101000000000000001000011;
		mem_i[65] = 32'b00011111100000000000000000000000;
		mem_i[66] = 32'b00101011111000000000000000000000;
		*/
		
		/*
		// Minloc 10
		mem_i[0] = 32'b00000000000000000000000000000000;
		mem_i[1] = 32'b00010111101000000010010101100000;
		mem_i[2] = 32'b00000111101111111111111011000011;
		mem_i[3] = 32'b00000111101111111111111111100011;
		mem_i[4] = 32'b00011011101111110000000000000000;
		mem_i[5] = 32'b00000111101111111111111111100011;
		mem_i[6] = 32'b00011011101111000000000000000000;
		mem_i[7] = 32'b00010011100111010000000000000000;
		mem_i[8] = 32'b00000111101111111111111111100011;
		mem_i[9] = 32'b00010001010111000000000000000000;
		mem_i[10] = 32'b00011101010000001111111111111111;
		mem_i[11] = 32'b00010101010000000000000000000000;
		mem_i[12] = 32'b00011011100010101111111111111111;
		mem_i[13] = 32'b00010001011111000000000000000000;
		mem_i[14] = 32'b00011101011000001111111111111111;
		mem_i[15] = 32'b00001101011000000000000101000111;
		mem_i[16] = 32'b00000111110000000000000000100011;
		mem_i[17] = 32'b00111100000000000000000000010001;
		mem_i[18] = 32'b00010101101000000010010101100000;
		mem_i[19] = 32'b00000101101010110000000000000010;
		mem_i[20] = 32'b00011101101000001111111111111111;
		mem_i[21] = 32'b00010111011000000000000000000000;
		mem_i[22] = 32'b01000011011000000000000000000000;
		mem_i[23] = 32'b00011111011000000000000000000000;
		mem_i[24] = 32'b00010001110110110000000000000000;
		mem_i[25] = 32'b00010001101011100000000000000000;
		mem_i[26] = 32'b00010111011000000010010101100000;
		mem_i[27] = 32'b00000111011010110000000000000010;
		mem_i[28] = 32'b00011011011011011111111111111111;
		mem_i[29] = 32'b00010011011010110000000000000000;
		mem_i[30] = 32'b00000111011000000000000000100011;
		mem_i[31] = 32'b00010001111110110000000000000000;
		mem_i[32] = 32'b00010001011011110000000000000000;
		mem_i[33] = 32'b00011011100010111111111111111111;
		mem_i[34] = 32'b00110100000000001111111111101010;
		mem_i[35] = 32'b00010110000000000010010101100000;
		mem_i[36] = 32'b00000110000111111111111111100011;
		mem_i[37] = 32'b00011011101010101111111111111111;
		mem_i[38] = 32'b00011011101010111111111111111110;
		mem_i[39] = 32'b00011011101011011111111111111101;
		mem_i[40] = 32'b00011011101100001111111111111100;
		mem_i[41] = 32'b00000111101111111111111110000011;
		mem_i[42] = 32'b00010111011000000000000101000000;
		mem_i[43] = 32'b00011011101110111111111111111011;
		mem_i[44] = 32'b00010111011000000000000000000000;
		mem_i[45] = 32'b00011011101110111111111111111100;
		mem_i[46] = 32'b00011011101100001111111111111101;
		mem_i[47] = 32'b00111000000000000000000000100000;
		mem_i[48] = 32'b00010010000111010000000000000000;
		mem_i[49] = 32'b00011110000000000000000000000000;
		mem_i[50] = 32'b00010001101111010000000000000000;
		mem_i[51] = 32'b00011101101000000000000000000001;
		mem_i[52] = 32'b00010001011111010000000000000000;
		mem_i[53] = 32'b00011101011000000000000000000010;
		mem_i[54] = 32'b00010001010111010000000000000000;
		mem_i[55] = 32'b00011101010000000000000000000011;
		mem_i[56] = 32'b00000111101000000000000010000011;
		mem_i[57] = 32'b00010010001110100000000000000000;
		mem_i[58] = 32'b00010010010111000000000000000000;
		mem_i[59] = 32'b00011110010000001111111111111111;
		mem_i[60] = 32'b00010110010000000000000000000000;
		mem_i[61] = 32'b00011011100100101111111111111111;
		mem_i[62] = 32'b00010010011111000000000000000000;
		mem_i[63] = 32'b00011110011000001111111111111111;
		mem_i[64] = 32'b00001110011000000000000101000111;
		mem_i[65] = 32'b00000111110000000000000000100011;
		mem_i[66] = 32'b00111100000000000000000000001100;
		mem_i[67] = 32'b00010110101000000010010101100000;
		mem_i[68] = 32'b00000110101100110000000000000010;
		mem_i[69] = 32'b00011110101000001111111111111111;
		mem_i[70] = 32'b00010111011000000000000000100000;
		mem_i[71] = 32'b00011011011101010000000000000000;
		mem_i[72] = 32'b01000111011000000000000000000000;
		mem_i[73] = 32'b00010011011100110000000000000000;
		mem_i[74] = 32'b00000111011000000000000000100011;
		mem_i[75] = 32'b00010010111110110000000000000000;
		mem_i[76] = 32'b00010010011101110000000000000000;
		mem_i[77] = 32'b00011011100100111111111111111111;
		mem_i[78] = 32'b00110100000000001111111111101111;
		mem_i[79] = 32'b11111100000000000000000000000000;
		mem_i[80] = 32'b00000111101111111111111111100011;
		mem_i[81] = 32'b00011011101111110000000000000000;
		mem_i[82] = 32'b00000111101111111111111111100011;
		mem_i[83] = 32'b00011011101111000000000000000000;
		mem_i[84] = 32'b00010011100111010000000000000000;
		mem_i[85] = 32'b00000111101111111111111111100011;
		mem_i[86] = 32'b00000111101111111111111111100011;
		mem_i[87] = 32'b00010010010111000000000000000000;
		mem_i[88] = 32'b00011110010000001111111111111110;
		mem_i[89] = 32'b00000111101111111111111111100011;
		mem_i[90] = 32'b00010010011111000000000000000000;
		mem_i[91] = 32'b00011110011000001111111111111101;
		mem_i[92] = 32'b00000111101111111111111111100011;
		mem_i[93] = 32'b00000111101111111111111111100011;
		mem_i[94] = 32'b00010010100111000000000000000000;
		mem_i[95] = 32'b00011110100000001111111111111100;
		mem_i[96] = 32'b00010010100100100000000000000000;
		mem_i[97] = 32'b00011011100101001111111111111100;
		mem_i[98] = 32'b00010010101111000000000000000000;
		mem_i[99] = 32'b00011110101000001111111111111100;
		mem_i[100] = 32'b00010010110111000000000000000000;
		mem_i[101] = 32'b00011110110000001111111111111101;
		mem_i[102] = 32'b00010011011101100000000000000000;
		mem_i[103] = 32'b00000111011000000000000000100100;
		mem_i[104] = 32'b00010010111110110000000000000000;
		mem_i[105] = 32'b00001110101101110000000000000001;
		mem_i[106] = 32'b00000111110000000000000000100011;
		mem_i[107] = 32'b00111100000000000000000001001100;
		mem_i[108] = 32'b00000111101111111111111111100011;
		mem_i[109] = 32'b00010011001111000000000000000000;
		mem_i[110] = 32'b00011111001000001111111111111011;
		mem_i[111] = 32'b00010000000111000000000000000000;
		mem_i[112] = 32'b00011100000000001111111111111111;
		mem_i[113] = 32'b00011011101000001111111111111111;
		mem_i[114] = 32'b00011011101100101111111111111110;
		mem_i[115] = 32'b00011011101100111111111111111101;
		mem_i[116] = 32'b00011011101101001111111111111100;
		mem_i[117] = 32'b00011011101101011111111111111011;
		mem_i[118] = 32'b00011011101101101111111111111010;
		mem_i[119] = 32'b00011011101110011111111111111001;
		mem_i[120] = 32'b00000111101111111111111100100011;
		mem_i[121] = 32'b00011011101101101111111111111011;
		mem_i[122] = 32'b00011011101101011111111111111100;
		mem_i[123] = 32'b00011011101000001111111111111101;
		mem_i[124] = 32'b00111000000000000000000001000001;
		mem_i[125] = 32'b00010011001111010000000000000000;
		mem_i[126] = 32'b00011111001000000000000000000000;
		mem_i[127] = 32'b00010010110111010000000000000000;
		mem_i[128] = 32'b00011110110000000000000000000001;
		mem_i[129] = 32'b00010010101111010000000000000000;
		mem_i[130] = 32'b00011110101000000000000000000010;
		mem_i[131] = 32'b00010010100111010000000000000000;
		mem_i[132] = 32'b00011110100000000000000000000011;
		mem_i[133] = 32'b00010010011111010000000000000000;
		mem_i[134] = 32'b00011110011000000000000000000100;
		mem_i[135] = 32'b00010010010111010000000000000000;
		mem_i[136] = 32'b00011110010000000000000000000101;
		mem_i[137] = 32'b00010000000111010000000000000000;
		mem_i[138] = 32'b00011100000000000000000000000110;
		mem_i[139] = 32'b00000111101000000000000011100011;
		mem_i[140] = 32'b00010000001110100000000000000000;
		mem_i[141] = 32'b00010011001000010000000000000000;
		mem_i[142] = 32'b00011011100110011111111111111011;
		mem_i[143] = 32'b00010000010111000000000000000000;
		mem_i[144] = 32'b00011100010000001111111111111010;
		mem_i[145] = 32'b00010000011111000000000000000000;
		mem_i[146] = 32'b00011100011000001111111111111011;
		mem_i[147] = 32'b00010000100111000000000000000000;
		mem_i[148] = 32'b00011100100000001111111111111111;
		mem_i[149] = 32'b00000100100000110000000000000010;
		mem_i[150] = 32'b00011100100000000000000000000000;
		mem_i[151] = 32'b00010000010001000000000000000000;
		mem_i[152] = 32'b00011011100000101111111111111010;
		mem_i[153] = 32'b00010000101111000000000000000000;
		mem_i[154] = 32'b00011100101000001111111111111111;
		mem_i[155] = 32'b00000100101000110000000000000010;
		mem_i[156] = 32'b00011100101000000000000000000000;
		mem_i[157] = 32'b00010000110111000000000000000000;
		mem_i[158] = 32'b00011100110000001111111111111100;
		mem_i[159] = 32'b00010000111111000000000000000000;
		mem_i[160] = 32'b00011100111000001111111111111111;
		mem_i[161] = 32'b00000100111001100000000000000010;
		mem_i[162] = 32'b00011100111000000000000000000000;
		mem_i[163] = 32'b00010000101001110000000000000000;
		mem_i[164] = 32'b00010011011111000000000000000000;
		mem_i[165] = 32'b00011111011000001111111111111111;
		mem_i[166] = 32'b00000111011000110000000000000010;
		mem_i[167] = 32'b00011011011001010000000000000000;
		mem_i[168] = 32'b00010001000111000000000000000000;
		mem_i[169] = 32'b00011101000000001111111111111111;
		mem_i[170] = 32'b00000101000001100000000000000010;
		mem_i[171] = 32'b00011101000000000000000000000000;
		mem_i[172] = 32'b00010001000000100000000000000000;
		mem_i[173] = 32'b00010011011111000000000000000000;
		mem_i[174] = 32'b00011111011000001111111111111111;
		mem_i[175] = 32'b00000111011001100000000000000010;
		mem_i[176] = 32'b00011011011010000000000000000000;
		mem_i[177] = 32'b00010011011001100000000000000000;
		mem_i[178] = 32'b00000111011000000000000000100011;
		mem_i[179] = 32'b00010001001110110000000000000000;
		mem_i[180] = 32'b00010000110010010000000000000000;
		mem_i[181] = 32'b00011011100001101111111111111100;
		mem_i[182] = 32'b00000111101000000000000000100011;
		mem_i[183] = 32'b00110100000000001111111110101010;
		mem_i[184] = 32'b00010011111111000000000000000000;
		mem_i[185] = 32'b00011111111000000000000000000001;
		mem_i[186] = 32'b00010011101111000000000000000000;
		mem_i[187] = 32'b00000111101000000000000001000011;
		mem_i[188] = 32'b00011111100000000000000000000000;
		mem_i[189] = 32'b00101011111000000000000000000000;
		mem_i[190] = 32'b00000111101111111111111111100011;
		mem_i[191] = 32'b00011011101111110000000000000000;
		mem_i[192] = 32'b00000111101111111111111111100011;
		mem_i[193] = 32'b00011011101111000000000000000000;
		mem_i[194] = 32'b00010011100111010000000000000000;
		mem_i[195] = 32'b00000111101111111111111111100011;
		mem_i[196] = 32'b00000111101111111111111111100011;
		mem_i[197] = 32'b00010000000111000000000000000000;
		mem_i[198] = 32'b00011100000000001111111111111110;
		mem_i[199] = 32'b00000111101111111111111111100011;
		mem_i[200] = 32'b00010000001111000000000000000000;
		mem_i[201] = 32'b00011100001000001111111111111101;
		mem_i[202] = 32'b00000111101111111111111111100011;
		mem_i[203] = 32'b00000111101111111111111111100011;
		mem_i[204] = 32'b00000111101111111111111111100011;
		mem_i[205] = 32'b00010000010111000000000000000000;
		mem_i[206] = 32'b00011100010000001111111111111010;
		mem_i[207] = 32'b00010000010000000000000000000000;
		mem_i[208] = 32'b00011011100000101111111111111010;
		mem_i[209] = 32'b00010000011111000000000000000000;
		mem_i[210] = 32'b00011100011000001111111111111011;
		mem_i[211] = 32'b00010000100111000000000000000000;
		mem_i[212] = 32'b00011100100000001111111111111111;
		mem_i[213] = 32'b00000100100000000000000000000010;
		mem_i[214] = 32'b00011100100000000000000000000000;
		mem_i[215] = 32'b00010000011001000000000000000000;
		mem_i[216] = 32'b00011011100000111111111111111011;
		mem_i[217] = 32'b00010000101111000000000000000000;
		mem_i[218] = 32'b00011100101000001111111111111100;
		mem_i[219] = 32'b00010011011000000000000000000000;
		mem_i[220] = 32'b00000111011000000000000000100011;
		mem_i[221] = 32'b00010000110110110000000000000000;
		mem_i[222] = 32'b00010000101001100000000000000000;
		mem_i[223] = 32'b00011011100001011111111111111100;
		mem_i[224] = 32'b00010000111111000000000000000000;
		mem_i[225] = 32'b00011100111000001111111111111100;
		mem_i[226] = 32'b00010001000111000000000000000000;
		mem_i[227] = 32'b00011101000000001111111111111101;
		mem_i[228] = 32'b00001100111010000000000000000001;
		mem_i[229] = 32'b00000111110000000000000000100011;
		mem_i[230] = 32'b00111100000000000000000000011100;
		mem_i[231] = 32'b00010001010111000000000000000000;
		mem_i[232] = 32'b00011101010000001111111111111111;
		mem_i[233] = 32'b00000101010001110000000000000010;
		mem_i[234] = 32'b00011101010000000000000000000000;
		mem_i[235] = 32'b00010001011111000000000000000000;
		mem_i[236] = 32'b00011101011000001111111111111011;
		mem_i[237] = 32'b00001101010010110000000000000001;
		mem_i[238] = 32'b00000111110000000000000000100011;
		mem_i[239] = 32'b00111100000000000000000000001011;
		mem_i[240] = 32'b00010001101111000000000000000000;
		mem_i[241] = 32'b00011101101000001111111111111111;
		mem_i[242] = 32'b00000101101001110000000000000010;
		mem_i[243] = 32'b00011101101000000000000000000000;
		mem_i[244] = 32'b00010001011011010000000000000000;
		mem_i[245] = 32'b00011011100010111111111111111011;
		mem_i[246] = 32'b00010001110111000000000000000000;
		mem_i[247] = 32'b00011101110000001111111111111010;
		mem_i[248] = 32'b00010001110001110000000000000000;
		mem_i[249] = 32'b00011011100011101111111111111010;
		mem_i[250] = 32'b00110100000000000000000000000000;
		mem_i[251] = 32'b00010001111111000000000000000000;
		mem_i[252] = 32'b00011101111000001111111111111100;
		mem_i[253] = 32'b00010011011011110000000000000000;
		mem_i[254] = 32'b00000111011000000000000000100011;
		mem_i[255] = 32'b00010010000110110000000000000000;
		mem_i[256] = 32'b00010001111100000000000000000000;
		mem_i[257] = 32'b00011011100011111111111111111100;
		mem_i[258] = 32'b00110100000000001111111111011101;
		mem_i[259] = 32'b00010010001111000000000000000000;
		mem_i[260] = 32'b00011110001000001111111111111010;
		mem_i[261] = 32'b00010011010100010000000000000000;
		mem_i[262] = 32'b00010011111111000000000000000000;
		mem_i[263] = 32'b00011111111000000000000000000001;
		mem_i[264] = 32'b00010011101111000000000000000000;
		mem_i[265] = 32'b00000111101000000000000001000011;
		mem_i[266] = 32'b00011111100000000000000000000000;
		mem_i[267] = 32'b00101011111000000000000000000000;
		*/
		
		/*
		// Minloc 5
		mem_i[0] = 32'b00000000000000000000000000000000;
		mem_i[1] = 32'b00010111101000000010010101100000;
		mem_i[2] = 32'b00000111101111111111111101100011;
		mem_i[3] = 32'b00000111101111111111111111100011;
		mem_i[4] = 32'b00011011101111110000000000000000;
		mem_i[5] = 32'b00000111101111111111111111100011;
		mem_i[6] = 32'b00011011101111000000000000000000;
		mem_i[7] = 32'b00010011100111010000000000000000;
		mem_i[8] = 32'b00000111101111111111111111100011;
		mem_i[9] = 32'b00010001010111000000000000000000;
		mem_i[10] = 32'b00011101010000001111111111111111;
		mem_i[11] = 32'b00010101010000000000000000000000;
		mem_i[12] = 32'b00011011100010101111111111111111;
		mem_i[13] = 32'b00010001011111000000000000000000;
		mem_i[14] = 32'b00011101011000001111111111111111;
		mem_i[15] = 32'b00001101011000000000000010100111;
		mem_i[16] = 32'b00000111110000000000000000100011;
		mem_i[17] = 32'b00111100000000000000000000010001;
		mem_i[18] = 32'b00010101101000000010010101100000;
		mem_i[19] = 32'b00000101101010110000000000000010;
		mem_i[20] = 32'b00011101101000001111111111111111;
		mem_i[21] = 32'b00010111011000000000000000000000;
		mem_i[22] = 32'b01000011011000000000000000000000;
		mem_i[23] = 32'b00011111011000000000000000000000;
		mem_i[24] = 32'b00010001110110110000000000000000;
		mem_i[25] = 32'b00010001101011100000000000000000;
		mem_i[26] = 32'b00010111011000000010010101100000;
		mem_i[27] = 32'b00000111011010110000000000000010;
		mem_i[28] = 32'b00011011011011011111111111111111;
		mem_i[29] = 32'b00010011011010110000000000000000;
		mem_i[30] = 32'b00000111011000000000000000100011;
		mem_i[31] = 32'b00010001111110110000000000000000;
		mem_i[32] = 32'b00010001011011110000000000000000;
		mem_i[33] = 32'b00011011100010111111111111111111;
		mem_i[34] = 32'b00110100000000001111111111101010;
		mem_i[35] = 32'b00010110000000000010010101100000;
		mem_i[36] = 32'b00000110000111111111111111100011;
		mem_i[37] = 32'b00011011101010101111111111111111;
		mem_i[38] = 32'b00011011101010111111111111111110;
		mem_i[39] = 32'b00011011101011011111111111111101;
		mem_i[40] = 32'b00011011101100001111111111111100;
		mem_i[41] = 32'b00000111101111111111111110000011;
		mem_i[42] = 32'b00010111011000000000000010100000;
		mem_i[43] = 32'b00011011101110111111111111111011;
		mem_i[44] = 32'b00010111011000000000000000000000;
		mem_i[45] = 32'b00011011101110111111111111111100;
		mem_i[46] = 32'b00011011101100001111111111111101;
		mem_i[47] = 32'b00111000000000000000000000100000;
		mem_i[48] = 32'b00010010000111010000000000000000;
		mem_i[49] = 32'b00011110000000000000000000000000;
		mem_i[50] = 32'b00010001101111010000000000000000;
		mem_i[51] = 32'b00011101101000000000000000000001;
		mem_i[52] = 32'b00010001011111010000000000000000;
		mem_i[53] = 32'b00011101011000000000000000000010;
		mem_i[54] = 32'b00010001010111010000000000000000;
		mem_i[55] = 32'b00011101010000000000000000000011;
		mem_i[56] = 32'b00000111101000000000000010000011;
		mem_i[57] = 32'b00010010001110100000000000000000;
		mem_i[58] = 32'b00010010010111000000000000000000;
		mem_i[59] = 32'b00011110010000001111111111111111;
		mem_i[60] = 32'b00010110010000000000000000000000;
		mem_i[61] = 32'b00011011100100101111111111111111;
		mem_i[62] = 32'b00010010011111000000000000000000;
		mem_i[63] = 32'b00011110011000001111111111111111;
		mem_i[64] = 32'b00001110011000000000000010100111;
		mem_i[65] = 32'b00000111110000000000000000100011;
		mem_i[66] = 32'b00111100000000000000000000001100;
		mem_i[67] = 32'b00010110101000000010010101100000;
		mem_i[68] = 32'b00000110101100110000000000000010;
		mem_i[69] = 32'b00011110101000001111111111111111;
		mem_i[70] = 32'b00010111011000000000000000100000;
		mem_i[71] = 32'b00011011011101010000000000000000;
		mem_i[72] = 32'b01000111011000000000000000000000;
		mem_i[73] = 32'b00010011011100110000000000000000;
		mem_i[74] = 32'b00000111011000000000000000100011;
		mem_i[75] = 32'b00010010111110110000000000000000;
		mem_i[76] = 32'b00010010011101110000000000000000;
		mem_i[77] = 32'b00011011100100111111111111111111;
		mem_i[78] = 32'b00110100000000001111111111101111;
		mem_i[79] = 32'b11111100000000000000000000000000;
		mem_i[80] = 32'b00000111101111111111111111100011;
		mem_i[81] = 32'b00011011101111110000000000000000;
		mem_i[82] = 32'b00000111101111111111111111100011;
		mem_i[83] = 32'b00011011101111000000000000000000;
		mem_i[84] = 32'b00010011100111010000000000000000;
		mem_i[85] = 32'b00000111101111111111111111100011;
		mem_i[86] = 32'b00000111101111111111111111100011;
		mem_i[87] = 32'b00010010010111000000000000000000;
		mem_i[88] = 32'b00011110010000001111111111111110;
		mem_i[89] = 32'b00000111101111111111111111100011;
		mem_i[90] = 32'b00010010011111000000000000000000;
		mem_i[91] = 32'b00011110011000001111111111111101;
		mem_i[92] = 32'b00000111101111111111111111100011;
		mem_i[93] = 32'b00000111101111111111111111100011;
		mem_i[94] = 32'b00010010100111000000000000000000;
		mem_i[95] = 32'b00011110100000001111111111111100;
		mem_i[96] = 32'b00010010100100100000000000000000;
		mem_i[97] = 32'b00011011100101001111111111111100;
		mem_i[98] = 32'b00010010101111000000000000000000;
		mem_i[99] = 32'b00011110101000001111111111111100;
		mem_i[100] = 32'b00010010110111000000000000000000;
		mem_i[101] = 32'b00011110110000001111111111111101;
		mem_i[102] = 32'b00010011011101100000000000000000;
		mem_i[103] = 32'b00000111011000000000000000100100;
		mem_i[104] = 32'b00010010111110110000000000000000;
		mem_i[105] = 32'b00001110101101110000000000000001;
		mem_i[106] = 32'b00000111110000000000000000100011;
		mem_i[107] = 32'b00111100000000000000000001001100;
		mem_i[108] = 32'b00000111101111111111111111100011;
		mem_i[109] = 32'b00010011001111000000000000000000;
		mem_i[110] = 32'b00011111001000001111111111111011;
		mem_i[111] = 32'b00010000000111000000000000000000;
		mem_i[112] = 32'b00011100000000001111111111111111;
		mem_i[113] = 32'b00011011101000001111111111111111;
		mem_i[114] = 32'b00011011101100101111111111111110;
		mem_i[115] = 32'b00011011101100111111111111111101;
		mem_i[116] = 32'b00011011101101001111111111111100;
		mem_i[117] = 32'b00011011101101011111111111111011;
		mem_i[118] = 32'b00011011101101101111111111111010;
		mem_i[119] = 32'b00011011101110011111111111111001;
		mem_i[120] = 32'b00000111101111111111111100100011;
		mem_i[121] = 32'b00011011101101101111111111111011;
		mem_i[122] = 32'b00011011101101011111111111111100;
		mem_i[123] = 32'b00011011101000001111111111111101;
		mem_i[124] = 32'b00111000000000000000000001000001;
		mem_i[125] = 32'b00010011001111010000000000000000;
		mem_i[126] = 32'b00011111001000000000000000000000;
		mem_i[127] = 32'b00010010110111010000000000000000;
		mem_i[128] = 32'b00011110110000000000000000000001;
		mem_i[129] = 32'b00010010101111010000000000000000;
		mem_i[130] = 32'b00011110101000000000000000000010;
		mem_i[131] = 32'b00010010100111010000000000000000;
		mem_i[132] = 32'b00011110100000000000000000000011;
		mem_i[133] = 32'b00010010011111010000000000000000;
		mem_i[134] = 32'b00011110011000000000000000000100;
		mem_i[135] = 32'b00010010010111010000000000000000;
		mem_i[136] = 32'b00011110010000000000000000000101;
		mem_i[137] = 32'b00010000000111010000000000000000;
		mem_i[138] = 32'b00011100000000000000000000000110;
		mem_i[139] = 32'b00000111101000000000000011100011;
		mem_i[140] = 32'b00010000001110100000000000000000;
		mem_i[141] = 32'b00010011001000010000000000000000;
		mem_i[142] = 32'b00011011100110011111111111111011;
		mem_i[143] = 32'b00010000010111000000000000000000;
		mem_i[144] = 32'b00011100010000001111111111111010;
		mem_i[145] = 32'b00010000011111000000000000000000;
		mem_i[146] = 32'b00011100011000001111111111111011;
		mem_i[147] = 32'b00010000100111000000000000000000;
		mem_i[148] = 32'b00011100100000001111111111111111;
		mem_i[149] = 32'b00000100100000110000000000000010;
		mem_i[150] = 32'b00011100100000000000000000000000;
		mem_i[151] = 32'b00010000010001000000000000000000;
		mem_i[152] = 32'b00011011100000101111111111111010;
		mem_i[153] = 32'b00010000101111000000000000000000;
		mem_i[154] = 32'b00011100101000001111111111111111;
		mem_i[155] = 32'b00000100101000110000000000000010;
		mem_i[156] = 32'b00011100101000000000000000000000;
		mem_i[157] = 32'b00010000110111000000000000000000;
		mem_i[158] = 32'b00011100110000001111111111111100;
		mem_i[159] = 32'b00010000111111000000000000000000;
		mem_i[160] = 32'b00011100111000001111111111111111;
		mem_i[161] = 32'b00000100111001100000000000000010;
		mem_i[162] = 32'b00011100111000000000000000000000;
		mem_i[163] = 32'b00010000101001110000000000000000;
		mem_i[164] = 32'b00010011011111000000000000000000;
		mem_i[165] = 32'b00011111011000001111111111111111;
		mem_i[166] = 32'b00000111011000110000000000000010;
		mem_i[167] = 32'b00011011011001010000000000000000;
		mem_i[168] = 32'b00010001000111000000000000000000;
		mem_i[169] = 32'b00011101000000001111111111111111;
		mem_i[170] = 32'b00000101000001100000000000000010;
		mem_i[171] = 32'b00011101000000000000000000000000;
		mem_i[172] = 32'b00010001000000100000000000000000;
		mem_i[173] = 32'b00010011011111000000000000000000;
		mem_i[174] = 32'b00011111011000001111111111111111;
		mem_i[175] = 32'b00000111011001100000000000000010;
		mem_i[176] = 32'b00011011011010000000000000000000;
		mem_i[177] = 32'b00010011011001100000000000000000;
		mem_i[178] = 32'b00000111011000000000000000100011;
		mem_i[179] = 32'b00010001001110110000000000000000;
		mem_i[180] = 32'b00010000110010010000000000000000;
		mem_i[181] = 32'b00011011100001101111111111111100;
		mem_i[182] = 32'b00000111101000000000000000100011;
		mem_i[183] = 32'b00110100000000001111111110101010;
		mem_i[184] = 32'b00010011111111000000000000000000;
		mem_i[185] = 32'b00011111111000000000000000000001;
		mem_i[186] = 32'b00010011101111000000000000000000;
		mem_i[187] = 32'b00000111101000000000000001000011;
		mem_i[188] = 32'b00011111100000000000000000000000;
		mem_i[189] = 32'b00101011111000000000000000000000;
		mem_i[190] = 32'b00000111101111111111111111100011;
		mem_i[191] = 32'b00011011101111110000000000000000;
		mem_i[192] = 32'b00000111101111111111111111100011;
		mem_i[193] = 32'b00011011101111000000000000000000;
		mem_i[194] = 32'b00010011100111010000000000000000;
		mem_i[195] = 32'b00000111101111111111111111100011;
		mem_i[196] = 32'b00000111101111111111111111100011;
		mem_i[197] = 32'b00010000000111000000000000000000;
		mem_i[198] = 32'b00011100000000001111111111111110;
		mem_i[199] = 32'b00000111101111111111111111100011;
		mem_i[200] = 32'b00010000001111000000000000000000;
		mem_i[201] = 32'b00011100001000001111111111111101;
		mem_i[202] = 32'b00000111101111111111111111100011;
		mem_i[203] = 32'b00000111101111111111111111100011;
		mem_i[204] = 32'b00000111101111111111111111100011;
		mem_i[205] = 32'b00010000010111000000000000000000;
		mem_i[206] = 32'b00011100010000001111111111111010;
		mem_i[207] = 32'b00010000010000000000000000000000;
		mem_i[208] = 32'b00011011100000101111111111111010;
		mem_i[209] = 32'b00010000011111000000000000000000;
		mem_i[210] = 32'b00011100011000001111111111111011;
		mem_i[211] = 32'b00010000100111000000000000000000;
		mem_i[212] = 32'b00011100100000001111111111111111;
		mem_i[213] = 32'b00000100100000000000000000000010;
		mem_i[214] = 32'b00011100100000000000000000000000;
		mem_i[215] = 32'b00010000011001000000000000000000;
		mem_i[216] = 32'b00011011100000111111111111111011;
		mem_i[217] = 32'b00010000101111000000000000000000;
		mem_i[218] = 32'b00011100101000001111111111111100;
		mem_i[219] = 32'b00010011011000000000000000000000;
		mem_i[220] = 32'b00000111011000000000000000100011;
		mem_i[221] = 32'b00010000110110110000000000000000;
		mem_i[222] = 32'b00010000101001100000000000000000;
		mem_i[223] = 32'b00011011100001011111111111111100;
		mem_i[224] = 32'b00010000111111000000000000000000;
		mem_i[225] = 32'b00011100111000001111111111111100;
		mem_i[226] = 32'b00010001000111000000000000000000;
		mem_i[227] = 32'b00011101000000001111111111111101;
		mem_i[228] = 32'b00001100111010000000000000000001;
		mem_i[229] = 32'b00000111110000000000000000100011;
		mem_i[230] = 32'b00111100000000000000000000011100;
		mem_i[231] = 32'b00010001010111000000000000000000;
		mem_i[232] = 32'b00011101010000001111111111111111;
		mem_i[233] = 32'b00000101010001110000000000000010;
		mem_i[234] = 32'b00011101010000000000000000000000;
		mem_i[235] = 32'b00010001011111000000000000000000;
		mem_i[236] = 32'b00011101011000001111111111111011;
		mem_i[237] = 32'b00001101010010110000000000000001;
		mem_i[238] = 32'b00000111110000000000000000100011;
		mem_i[239] = 32'b00111100000000000000000000001011;
		mem_i[240] = 32'b00010001101111000000000000000000;
		mem_i[241] = 32'b00011101101000001111111111111111;
		mem_i[242] = 32'b00000101101001110000000000000010;
		mem_i[243] = 32'b00011101101000000000000000000000;
		mem_i[244] = 32'b00010001011011010000000000000000;
		mem_i[245] = 32'b00011011100010111111111111111011;
		mem_i[246] = 32'b00010001110111000000000000000000;
		mem_i[247] = 32'b00011101110000001111111111111010;
		mem_i[248] = 32'b00010001110001110000000000000000;
		mem_i[249] = 32'b00011011100011101111111111111010;
		mem_i[250] = 32'b00110100000000000000000000000000;
		mem_i[251] = 32'b00010001111111000000000000000000;
		mem_i[252] = 32'b00011101111000001111111111111100;
		mem_i[253] = 32'b00010011011011110000000000000000;
		mem_i[254] = 32'b00000111011000000000000000100011;
		mem_i[255] = 32'b00010010000110110000000000000000;
		mem_i[256] = 32'b00010001111100000000000000000000;
		mem_i[257] = 32'b00011011100011111111111111111100;
		mem_i[258] = 32'b00110100000000001111111111011101;
		mem_i[259] = 32'b00010010001111000000000000000000;
		mem_i[260] = 32'b00011110001000001111111111111010;
		mem_i[261] = 32'b00010011010100010000000000000000;
		mem_i[262] = 32'b00010011111111000000000000000000;
		mem_i[263] = 32'b00011111111000000000000000000001;
		mem_i[264] = 32'b00010011101111000000000000000000;
		mem_i[265] = 32'b00000111101000000000000001000011;
		mem_i[266] = 32'b00011111100000000000000000000000;
		mem_i[267] = 32'b00101011111000000000000000000000;
		*/
	
		// Minloc 3
		/*
		mem_i[0] = 32'b00000000000000000000000000000000;
		mem_i[1] = 32'b00010111101000000010010101100000;
		mem_i[2] = 32'b00000111101111111111111110100011;
		mem_i[3] = 32'b00000111101111111111111111100011;
		mem_i[4] = 32'b00011011101111110000000000000000;
		mem_i[5] = 32'b00000111101111111111111111100011;
		mem_i[6] = 32'b00011011101111000000000000000000;
		mem_i[7] = 32'b00010011100111010000000000000000;
		mem_i[8] = 32'b00000111101111111111111111100011;
		mem_i[9] = 32'b00010001010111000000000000000000;
		mem_i[10] = 32'b00011101010000001111111111111111;
		mem_i[11] = 32'b00010101010000000000000000000000;
		mem_i[12] = 32'b00011011100010101111111111111111;
		mem_i[13] = 32'b00010001011111000000000000000000;
		mem_i[14] = 32'b00011101011000001111111111111111;
		mem_i[15] = 32'b00001101011000000000000001100111;
		mem_i[16] = 32'b00000111110000000000000000100011;
		mem_i[17] = 32'b00111100000000000000000000010001;
		mem_i[18] = 32'b00010101101000000010010101100000;
		mem_i[19] = 32'b00000101101010110000000000000010;
		mem_i[20] = 32'b00011101101000001111111111111111;
		mem_i[21] = 32'b00010111011000000000000000000000;
		mem_i[22] = 32'b01000011011000000000000000000000;
		mem_i[23] = 32'b00011111011000000000000000000000;
		mem_i[24] = 32'b00010001110110110000000000000000;
		mem_i[25] = 32'b00010001101011100000000000000000;
		mem_i[26] = 32'b00010111011000000010010101100000;
		mem_i[27] = 32'b00000111011010110000000000000010;
		mem_i[28] = 32'b00011011011011011111111111111111;
		mem_i[29] = 32'b00010011011010110000000000000000;
		mem_i[30] = 32'b00000111011000000000000000100011;
		mem_i[31] = 32'b00010001111110110000000000000000;
		mem_i[32] = 32'b00010001011011110000000000000000;
		mem_i[33] = 32'b00011011100010111111111111111111;
		mem_i[34] = 32'b00110100000000001111111111101010;
		mem_i[35] = 32'b00010110000000000010010101100000;
		mem_i[36] = 32'b00000110000111111111111111100011;
		mem_i[37] = 32'b00011011101010101111111111111111;
		mem_i[38] = 32'b00011011101010111111111111111110;
		mem_i[39] = 32'b00011011101011011111111111111101;
		mem_i[40] = 32'b00011011101100001111111111111100;
		mem_i[41] = 32'b00000111101111111111111110000011;
		mem_i[42] = 32'b00010111011000000000000001100000;
		mem_i[43] = 32'b00011011101110111111111111111011;
		mem_i[44] = 32'b00010111011000000000000000000000;
		mem_i[45] = 32'b00011011101110111111111111111100;
		mem_i[46] = 32'b00011011101100001111111111111101;
		mem_i[47] = 32'b00111000000000000000000000100000;
		mem_i[48] = 32'b00010010000111010000000000000000;
		mem_i[49] = 32'b00011110000000000000000000000000;
		mem_i[50] = 32'b00010001101111010000000000000000;
		mem_i[51] = 32'b00011101101000000000000000000001;
		mem_i[52] = 32'b00010001011111010000000000000000;
		mem_i[53] = 32'b00011101011000000000000000000010;
		mem_i[54] = 32'b00010001010111010000000000000000;
		mem_i[55] = 32'b00011101010000000000000000000011;
		mem_i[56] = 32'b00000111101000000000000010000011;
		mem_i[57] = 32'b00010010001110100000000000000000;
		mem_i[58] = 32'b00010010010111000000000000000000;
		mem_i[59] = 32'b00011110010000001111111111111111;
		mem_i[60] = 32'b00010110010000000000000000000000;
		mem_i[61] = 32'b00011011100100101111111111111111;
		mem_i[62] = 32'b00010010011111000000000000000000;
		mem_i[63] = 32'b00011110011000001111111111111111;
		mem_i[64] = 32'b00001110011000000000000001100111;
		mem_i[65] = 32'b00000111110000000000000000100011;
		mem_i[66] = 32'b00111100000000000000000000001100;
		mem_i[67] = 32'b00010110101000000010010101100000;
		mem_i[68] = 32'b00000110101100110000000000000010;
		mem_i[69] = 32'b00011110101000001111111111111111;
		mem_i[70] = 32'b00010111011000000000000000100000;
		mem_i[71] = 32'b00011011011101010000000000000000;
		mem_i[72] = 32'b01000111011000000000000000000000;
		mem_i[73] = 32'b00010011011100110000000000000000;
		mem_i[74] = 32'b00000111011000000000000000100011;
		mem_i[75] = 32'b00010010111110110000000000000000;
		mem_i[76] = 32'b00010010011101110000000000000000;
		mem_i[77] = 32'b00011011100100111111111111111111;
		mem_i[78] = 32'b00110100000000001111111111101111;
		mem_i[79] = 32'b11111100000000000000000000000000;
		mem_i[80] = 32'b00000111101111111111111111100011;
		mem_i[81] = 32'b00011011101111110000000000000000;
		mem_i[82] = 32'b00000111101111111111111111100011;
		mem_i[83] = 32'b00011011101111000000000000000000;
		mem_i[84] = 32'b00010011100111010000000000000000;
		mem_i[85] = 32'b00000111101111111111111111100011;
		mem_i[86] = 32'b00000111101111111111111111100011;
		mem_i[87] = 32'b00010010010111000000000000000000;
		mem_i[88] = 32'b00011110010000001111111111111110;
		mem_i[89] = 32'b00000111101111111111111111100011;
		mem_i[90] = 32'b00010010011111000000000000000000;
		mem_i[91] = 32'b00011110011000001111111111111101;
		mem_i[92] = 32'b00000111101111111111111111100011;
		mem_i[93] = 32'b00000111101111111111111111100011;
		mem_i[94] = 32'b00010010100111000000000000000000;
		mem_i[95] = 32'b00011110100000001111111111111100;
		mem_i[96] = 32'b00010010100100100000000000000000;
		mem_i[97] = 32'b00011011100101001111111111111100;
		mem_i[98] = 32'b00010010101111000000000000000000;
		mem_i[99] = 32'b00011110101000001111111111111100;
		mem_i[100] = 32'b00010010110111000000000000000000;
		mem_i[101] = 32'b00011110110000001111111111111101;
		mem_i[102] = 32'b00010011011101100000000000000000;
		mem_i[103] = 32'b00000111011000000000000000100100;
		mem_i[104] = 32'b00010010111110110000000000000000;
		mem_i[105] = 32'b00001110101101110000000000000001;
		mem_i[106] = 32'b00000111110000000000000000100011;
		mem_i[107] = 32'b00111100000000000000000001001100;
		mem_i[108] = 32'b00000111101111111111111111100011;
		mem_i[109] = 32'b00010011001111000000000000000000;
		mem_i[110] = 32'b00011111001000001111111111111011;
		mem_i[111] = 32'b00010000000111000000000000000000;
		mem_i[112] = 32'b00011100000000001111111111111111;
		mem_i[113] = 32'b00011011101000001111111111111111;
		mem_i[114] = 32'b00011011101100101111111111111110;
		mem_i[115] = 32'b00011011101100111111111111111101;
		mem_i[116] = 32'b00011011101101001111111111111100;
		mem_i[117] = 32'b00011011101101011111111111111011;
		mem_i[118] = 32'b00011011101101101111111111111010;
		mem_i[119] = 32'b00011011101110011111111111111001;
		mem_i[120] = 32'b00000111101111111111111100100011;
		mem_i[121] = 32'b00011011101101101111111111111011;
		mem_i[122] = 32'b00011011101101011111111111111100;
		mem_i[123] = 32'b00011011101000001111111111111101;
		mem_i[124] = 32'b00111000000000000000000001000001;
		mem_i[125] = 32'b00010011001111010000000000000000;
		mem_i[126] = 32'b00011111001000000000000000000000;
		mem_i[127] = 32'b00010010110111010000000000000000;
		mem_i[128] = 32'b00011110110000000000000000000001;
		mem_i[129] = 32'b00010010101111010000000000000000;
		mem_i[130] = 32'b00011110101000000000000000000010;
		mem_i[131] = 32'b00010010100111010000000000000000;
		mem_i[132] = 32'b00011110100000000000000000000011;
		mem_i[133] = 32'b00010010011111010000000000000000;
		mem_i[134] = 32'b00011110011000000000000000000100;
		mem_i[135] = 32'b00010010010111010000000000000000;
		mem_i[136] = 32'b00011110010000000000000000000101;
		mem_i[137] = 32'b00010000000111010000000000000000;
		mem_i[138] = 32'b00011100000000000000000000000110;
		mem_i[139] = 32'b00000111101000000000000011100011;
		mem_i[140] = 32'b00010000001110100000000000000000;
		mem_i[141] = 32'b00010011001000010000000000000000;
		mem_i[142] = 32'b00011011100110011111111111111011;
		mem_i[143] = 32'b00010000010111000000000000000000;
		mem_i[144] = 32'b00011100010000001111111111111010;
		mem_i[145] = 32'b00010000011111000000000000000000;
		mem_i[146] = 32'b00011100011000001111111111111011;
		mem_i[147] = 32'b00010000100111000000000000000000;
		mem_i[148] = 32'b00011100100000001111111111111111;
		mem_i[149] = 32'b00000100100000110000000000000010;
		mem_i[150] = 32'b00011100100000000000000000000000;
		mem_i[151] = 32'b00010000010001000000000000000000;
		mem_i[152] = 32'b00011011100000101111111111111010;
		mem_i[153] = 32'b00010000101111000000000000000000;
		mem_i[154] = 32'b00011100101000001111111111111111;
		mem_i[155] = 32'b00000100101000110000000000000010;
		mem_i[156] = 32'b00011100101000000000000000000000;
		mem_i[157] = 32'b00010000110111000000000000000000;
		mem_i[158] = 32'b00011100110000001111111111111100;
		mem_i[159] = 32'b00010000111111000000000000000000;
		mem_i[160] = 32'b00011100111000001111111111111111;
		mem_i[161] = 32'b00000100111001100000000000000010;
		mem_i[162] = 32'b00011100111000000000000000000000;
		mem_i[163] = 32'b00010000101001110000000000000000;
		mem_i[164] = 32'b00010011011111000000000000000000;
		mem_i[165] = 32'b00011111011000001111111111111111;
		mem_i[166] = 32'b00000111011000110000000000000010;
		mem_i[167] = 32'b00011011011001010000000000000000;
		mem_i[168] = 32'b00010001000111000000000000000000;
		mem_i[169] = 32'b00011101000000001111111111111111;
		mem_i[170] = 32'b00000101000001100000000000000010;
		mem_i[171] = 32'b00011101000000000000000000000000;
		mem_i[172] = 32'b00010001000000100000000000000000;
		mem_i[173] = 32'b00010011011111000000000000000000;
		mem_i[174] = 32'b00011111011000001111111111111111;
		mem_i[175] = 32'b00000111011001100000000000000010;
		mem_i[176] = 32'b00011011011010000000000000000000;
		mem_i[177] = 32'b00010011011001100000000000000000;
		mem_i[178] = 32'b00000111011000000000000000100011;
		mem_i[179] = 32'b00010001001110110000000000000000;
		mem_i[180] = 32'b00010000110010010000000000000000;
		mem_i[181] = 32'b00011011100001101111111111111100;
		mem_i[182] = 32'b00000111101000000000000000100011;
		mem_i[183] = 32'b00110100000000001111111110101010;
		mem_i[184] = 32'b00010011111111000000000000000000;
		mem_i[185] = 32'b00011111111000000000000000000001;
		mem_i[186] = 32'b00010011101111000000000000000000;
		mem_i[187] = 32'b00000111101000000000000001000011;
		mem_i[188] = 32'b00011111100000000000000000000000;
		mem_i[189] = 32'b00101011111000000000000000000000;
		mem_i[190] = 32'b00000111101111111111111111100011;
		mem_i[191] = 32'b00011011101111110000000000000000;
		mem_i[192] = 32'b00000111101111111111111111100011;
		mem_i[193] = 32'b00011011101111000000000000000000;
		mem_i[194] = 32'b00010011100111010000000000000000;
		mem_i[195] = 32'b00000111101111111111111111100011;
		mem_i[196] = 32'b00000111101111111111111111100011;
		mem_i[197] = 32'b00010000000111000000000000000000;
		mem_i[198] = 32'b00011100000000001111111111111110;
		mem_i[199] = 32'b00000111101111111111111111100011;
		mem_i[200] = 32'b00010000001111000000000000000000;
		mem_i[201] = 32'b00011100001000001111111111111101;
		mem_i[202] = 32'b00000111101111111111111111100011;
		mem_i[203] = 32'b00000111101111111111111111100011;
		mem_i[204] = 32'b00000111101111111111111111100011;
		mem_i[205] = 32'b00010000010111000000000000000000;
		mem_i[206] = 32'b00011100010000001111111111111010;
		mem_i[207] = 32'b00010000010000000000000000000000;
		mem_i[208] = 32'b00011011100000101111111111111010;
		mem_i[209] = 32'b00010000011111000000000000000000;
		mem_i[210] = 32'b00011100011000001111111111111011;
		mem_i[211] = 32'b00010000100111000000000000000000;
		mem_i[212] = 32'b00011100100000001111111111111111;
		mem_i[213] = 32'b00000100100000000000000000000010;
		mem_i[214] = 32'b00011100100000000000000000000000;
		mem_i[215] = 32'b00010000011001000000000000000000;
		mem_i[216] = 32'b00011011100000111111111111111011;
		mem_i[217] = 32'b00010000101111000000000000000000;
		mem_i[218] = 32'b00011100101000001111111111111100;
		mem_i[219] = 32'b00010011011000000000000000000000;
		mem_i[220] = 32'b00000111011000000000000000100011;
		mem_i[221] = 32'b00010000110110110000000000000000;
		mem_i[222] = 32'b00010000101001100000000000000000;
		mem_i[223] = 32'b00011011100001011111111111111100;
		mem_i[224] = 32'b00010000111111000000000000000000;
		mem_i[225] = 32'b00011100111000001111111111111100;
		mem_i[226] = 32'b00010001000111000000000000000000;
		mem_i[227] = 32'b00011101000000001111111111111101;
		mem_i[228] = 32'b00001100111010000000000000000001;
		mem_i[229] = 32'b00000111110000000000000000100011;
		mem_i[230] = 32'b00111100000000000000000000011100;
		mem_i[231] = 32'b00010001010111000000000000000000;
		mem_i[232] = 32'b00011101010000001111111111111111;
		mem_i[233] = 32'b00000101010001110000000000000010;
		mem_i[234] = 32'b00011101010000000000000000000000;
		mem_i[235] = 32'b00010001011111000000000000000000;
		mem_i[236] = 32'b00011101011000001111111111111011;
		mem_i[237] = 32'b00001101010010110000000000000001;
		mem_i[238] = 32'b00000111110000000000000000100011;
		mem_i[239] = 32'b00111100000000000000000000001011;
		mem_i[240] = 32'b00010001101111000000000000000000;
		mem_i[241] = 32'b00011101101000001111111111111111;
		mem_i[242] = 32'b00000101101001110000000000000010;
		mem_i[243] = 32'b00011101101000000000000000000000;
		mem_i[244] = 32'b00010001011011010000000000000000;
		mem_i[245] = 32'b00011011100010111111111111111011;
		mem_i[246] = 32'b00010001110111000000000000000000;
		mem_i[247] = 32'b00011101110000001111111111111010;
		mem_i[248] = 32'b00010001110001110000000000000000;
		mem_i[249] = 32'b00011011100011101111111111111010;
		mem_i[250] = 32'b00110100000000000000000000000000;
		mem_i[251] = 32'b00010001111111000000000000000000;
		mem_i[252] = 32'b00011101111000001111111111111100;
		mem_i[253] = 32'b00010011011011110000000000000000;
		mem_i[254] = 32'b00000111011000000000000000100011;
		mem_i[255] = 32'b00010010000110110000000000000000;
		mem_i[256] = 32'b00010001111100000000000000000000;
		mem_i[257] = 32'b00011011100011111111111111111100;
		mem_i[258] = 32'b00110100000000001111111111011101;
		mem_i[259] = 32'b00010010001111000000000000000000;
		mem_i[260] = 32'b00011110001000001111111111111010;
		mem_i[261] = 32'b00010011010100010000000000000000;
		mem_i[262] = 32'b00010011111111000000000000000000;
		mem_i[263] = 32'b00011111111000000000000000000001;
		mem_i[264] = 32'b00010011101111000000000000000000;
		mem_i[265] = 32'b00000111101000000000000001000011;
		mem_i[266] = 32'b00011111100000000000000000000000;
		mem_i[267] = 32'b00101011111000000000000000000000;
		*/


		/*
		// Fibonacci
		mem_i[0 ] = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;	// START
		mem_i[1 ] = 32'b00010100000000000000000000000000;
		mem_i[2 ] = 32'b01000000000000000000000000000000;
		mem_i[3 ] = 32'b00011100000000000000000000000000;
		mem_i[4 ] = 32'b00111000000000000000000000000101;	//bal
		mem_i[5 ] = 32'b00010000001011010000000000000000;
		mem_i[6 ] = 32'b00010100000000000000000000000000;
		mem_i[7 ] = 32'b00011000000000010000000000000000;
		mem_i[8 ] = 32'b01000100000000000000000000000000;
		mem_i[9 ] = 32'b11111100000000000000000000000000;	// STOP
		mem_i[10] = 32'b00010001010000000000000000000000;
		mem_i[11] = 32'b00010101011000000000000000000000;
		mem_i[12] = 32'b00010101100000000000000000100000;
		mem_i[13] = 32'b00010101101000000000000000100000;
		mem_i[14] = 32'b00001101010000000000000001001011;
		mem_i[15] = 32'b00110011111000000000000000000000;
		mem_i[16] = 32'b00000000000000000000000000000000;	// NOP
		mem_i[17] = 32'b00000101010000000000000001000100;
		mem_i[18] = 32'b00001101011010100000000000000110;
		mem_i[19] = 32'b00111100000000000000000000000101;	// branch afterfor
		mem_i[20] = 32'b00010001110011010000000000000000;	// mv r14, r13
		mem_i[21] = 32'b00000101101011000000000000000001;
		mem_i[22] = 32'b00010001100011100000000000000000;
		mem_i[23] = 32'b00000101011000000000000000100011;	// addi
		mem_i[24] = 32'b00110100000000001111111111111001;	// branch for
		mem_i[25] = 32'b00110011111000000000000000000000;	// jc 
		//mem_i[26] = 32'b;											// END
		*/
	
		/**/
		
	end
	
	assign ID = mem_i[I];   // Repassa dado do endereco I
	
endmodule
